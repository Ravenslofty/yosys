module \$_DFF_P_ (input D, C, output Q);
    wire _TECHMAP_REMOVEINIT_Q_ = 1;
    dff _TECHMAP_REPLACE_ (.Q(Q), .D(D), .CLK(C));
endmodule
